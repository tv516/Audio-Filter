-- nios_system.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity nios_system is
	port (
		AUD_ADCDAT_to_the_audio_0   : in    std_logic                     := '0';             --     audio.ADCDAT
		AUD_ADCLRCK_to_the_audio_0  : in    std_logic                     := '0';             --          .ADCLRCK
		AUD_BCLK_to_the_audio_0     : in    std_logic                     := '0';             --          .BCLK
		AUD_DACDAT_from_the_audio_0 : out   std_logic;                                        --          .DACDAT
		AUD_DACLRCK_to_the_audio_0  : in    std_logic                     := '0';             --          .DACLRCK
		clk_clk                     : in    std_logic                     := '0';             --       clk.clk
		i2c_SDAT                    : inout std_logic                     := '0';             --       i2c.SDAT
		i2c_SCLK                    : out   std_logic;                                        --          .SCLK
		pin_export                  : out   std_logic;                                        --       pin.export
		reset_reset                 : in    std_logic                     := '0';             --     reset.reset
		sdram_addr                  : out   std_logic_vector(12 downto 0);                    --     sdram.addr
		sdram_ba                    : out   std_logic_vector(1 downto 0);                     --          .ba
		sdram_cas_n                 : out   std_logic;                                        --          .cas_n
		sdram_cke                   : out   std_logic;                                        --          .cke
		sdram_cs_n                  : out   std_logic;                                        --          .cs_n
		sdram_dq                    : inout std_logic_vector(15 downto 0) := (others => '0'); --          .dq
		sdram_dqm                   : out   std_logic_vector(1 downto 0);                     --          .dqm
		sdram_ras_n                 : out   std_logic;                                        --          .ras_n
		sdram_we_n                  : out   std_logic;                                        --          .we_n
		sdram_clk_clk               : out   std_logic;                                        -- sdram_clk.clk
		sw_export                   : in    std_logic_vector(7 downto 0)  := (others => '0')  --        sw.export
	);
end entity nios_system;

architecture rtl of nios_system is
	component nios_system_audio_0 is
		port (
			clk         : in  std_logic                     := 'X';             -- clk
			reset       : in  std_logic                     := 'X';             -- reset
			address     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			chipselect  : in  std_logic                     := 'X';             -- chipselect
			read        : in  std_logic                     := 'X';             -- read
			write       : in  std_logic                     := 'X';             -- write
			writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			irq         : out std_logic;                                        -- irq
			AUD_ADCDAT  : in  std_logic                     := 'X';             -- export
			AUD_ADCLRCK : in  std_logic                     := 'X';             -- export
			AUD_BCLK    : in  std_logic                     := 'X';             -- export
			AUD_DACDAT  : out std_logic;                                        -- export
			AUD_DACLRCK : in  std_logic                     := 'X'              -- export
		);
	end component nios_system_audio_0;

	component nios_system_audio_and_video_config_0 is
		port (
			clk         : in    std_logic                     := 'X';             -- clk
			reset       : in    std_logic                     := 'X';             -- reset
			address     : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			byteenable  : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			read        : in    std_logic                     := 'X';             -- read
			write       : in    std_logic                     := 'X';             -- write
			writedata   : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			readdata    : out   std_logic_vector(31 downto 0);                    -- readdata
			waitrequest : out   std_logic;                                        -- waitrequest
			I2C_SDAT    : inout std_logic                     := 'X';             -- export
			I2C_SCLK    : out   std_logic                                         -- export
		);
	end component nios_system_audio_and_video_config_0;

	component nios_system_jtag_uart_0 is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component nios_system_jtag_uart_0;

	component nios_system_new_sdram_controller_0 is
		port (
			clk            : in    std_logic                     := 'X';             -- clk
			reset_n        : in    std_logic                     := 'X';             -- reset_n
			az_addr        : in    std_logic_vector(24 downto 0) := (others => 'X'); -- address
			az_be_n        : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable_n
			az_cs          : in    std_logic                     := 'X';             -- chipselect
			az_data        : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			az_rd_n        : in    std_logic                     := 'X';             -- read_n
			az_wr_n        : in    std_logic                     := 'X';             -- write_n
			za_data        : out   std_logic_vector(15 downto 0);                    -- readdata
			za_valid       : out   std_logic;                                        -- readdatavalid
			za_waitrequest : out   std_logic;                                        -- waitrequest
			zs_addr        : out   std_logic_vector(12 downto 0);                    -- export
			zs_ba          : out   std_logic_vector(1 downto 0);                     -- export
			zs_cas_n       : out   std_logic;                                        -- export
			zs_cke         : out   std_logic;                                        -- export
			zs_cs_n        : out   std_logic;                                        -- export
			zs_dq          : inout std_logic_vector(15 downto 0) := (others => 'X'); -- export
			zs_dqm         : out   std_logic_vector(1 downto 0);                     -- export
			zs_ras_n       : out   std_logic;                                        -- export
			zs_we_n        : out   std_logic                                         -- export
		);
	end component nios_system_new_sdram_controller_0;

	component nios_system_nios2_gen2_0 is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(26 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(26 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component nios_system_nios2_gen2_0;

	component nios_system_onchip_memory2_1 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(13 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			freeze     : in  std_logic                     := 'X'              -- freeze
		);
	end component nios_system_onchip_memory2_1;

	component nios_system_pin is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic                                         -- export
		);
	end component nios_system_pin;

	component nios_system_pio_0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_port    : in  std_logic_vector(7 downto 0)  := (others => 'X')  -- export
		);
	end component nios_system_pio_0;

	component nios_system_sys_sdram_pll_0 is
		port (
			ref_clk_clk        : in  std_logic := 'X'; -- clk
			ref_reset_reset    : in  std_logic := 'X'; -- reset
			sys_clk_clk        : out std_logic;        -- clk
			sdram_clk_clk      : out std_logic;        -- clk
			reset_source_reset : out std_logic         -- reset
		);
	end component nios_system_sys_sdram_pll_0;

	component nios_system_sysid is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component nios_system_sysid;

	component nios_system_timer_0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component nios_system_timer_0;

	component nios_system_mm_interconnect_0 is
		port (
			sys_sdram_pll_0_sys_clk_clk                                 : in  std_logic                     := 'X';             -- clk
			nios2_gen2_0_reset_reset_bridge_in_reset_reset              : in  std_logic                     := 'X';             -- reset
			nios2_gen2_0_data_master_address                            : in  std_logic_vector(26 downto 0) := (others => 'X'); -- address
			nios2_gen2_0_data_master_waitrequest                        : out std_logic;                                        -- waitrequest
			nios2_gen2_0_data_master_byteenable                         : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			nios2_gen2_0_data_master_read                               : in  std_logic                     := 'X';             -- read
			nios2_gen2_0_data_master_readdata                           : out std_logic_vector(31 downto 0);                    -- readdata
			nios2_gen2_0_data_master_write                              : in  std_logic                     := 'X';             -- write
			nios2_gen2_0_data_master_writedata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			nios2_gen2_0_data_master_debugaccess                        : in  std_logic                     := 'X';             -- debugaccess
			nios2_gen2_0_instruction_master_address                     : in  std_logic_vector(26 downto 0) := (others => 'X'); -- address
			nios2_gen2_0_instruction_master_waitrequest                 : out std_logic;                                        -- waitrequest
			nios2_gen2_0_instruction_master_read                        : in  std_logic                     := 'X';             -- read
			nios2_gen2_0_instruction_master_readdata                    : out std_logic_vector(31 downto 0);                    -- readdata
			audio_0_avalon_audio_slave_address                          : out std_logic_vector(1 downto 0);                     -- address
			audio_0_avalon_audio_slave_write                            : out std_logic;                                        -- write
			audio_0_avalon_audio_slave_read                             : out std_logic;                                        -- read
			audio_0_avalon_audio_slave_readdata                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			audio_0_avalon_audio_slave_writedata                        : out std_logic_vector(31 downto 0);                    -- writedata
			audio_0_avalon_audio_slave_chipselect                       : out std_logic;                                        -- chipselect
			audio_and_video_config_0_avalon_av_config_slave_address     : out std_logic_vector(1 downto 0);                     -- address
			audio_and_video_config_0_avalon_av_config_slave_write       : out std_logic;                                        -- write
			audio_and_video_config_0_avalon_av_config_slave_read        : out std_logic;                                        -- read
			audio_and_video_config_0_avalon_av_config_slave_readdata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			audio_and_video_config_0_avalon_av_config_slave_writedata   : out std_logic_vector(31 downto 0);                    -- writedata
			audio_and_video_config_0_avalon_av_config_slave_byteenable  : out std_logic_vector(3 downto 0);                     -- byteenable
			audio_and_video_config_0_avalon_av_config_slave_waitrequest : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_0_avalon_jtag_slave_address                       : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart_0_avalon_jtag_slave_write                         : out std_logic;                                        -- write
			jtag_uart_0_avalon_jtag_slave_read                          : out std_logic;                                        -- read
			jtag_uart_0_avalon_jtag_slave_readdata                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_0_avalon_jtag_slave_writedata                     : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_0_avalon_jtag_slave_waitrequest                   : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_0_avalon_jtag_slave_chipselect                    : out std_logic;                                        -- chipselect
			new_sdram_controller_0_s1_address                           : out std_logic_vector(24 downto 0);                    -- address
			new_sdram_controller_0_s1_write                             : out std_logic;                                        -- write
			new_sdram_controller_0_s1_read                              : out std_logic;                                        -- read
			new_sdram_controller_0_s1_readdata                          : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			new_sdram_controller_0_s1_writedata                         : out std_logic_vector(15 downto 0);                    -- writedata
			new_sdram_controller_0_s1_byteenable                        : out std_logic_vector(1 downto 0);                     -- byteenable
			new_sdram_controller_0_s1_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			new_sdram_controller_0_s1_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			new_sdram_controller_0_s1_chipselect                        : out std_logic;                                        -- chipselect
			nios2_gen2_0_debug_mem_slave_address                        : out std_logic_vector(8 downto 0);                     -- address
			nios2_gen2_0_debug_mem_slave_write                          : out std_logic;                                        -- write
			nios2_gen2_0_debug_mem_slave_read                           : out std_logic;                                        -- read
			nios2_gen2_0_debug_mem_slave_readdata                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nios2_gen2_0_debug_mem_slave_writedata                      : out std_logic_vector(31 downto 0);                    -- writedata
			nios2_gen2_0_debug_mem_slave_byteenable                     : out std_logic_vector(3 downto 0);                     -- byteenable
			nios2_gen2_0_debug_mem_slave_waitrequest                    : in  std_logic                     := 'X';             -- waitrequest
			nios2_gen2_0_debug_mem_slave_debugaccess                    : out std_logic;                                        -- debugaccess
			onchip_memory2_1_s1_address                                 : out std_logic_vector(13 downto 0);                    -- address
			onchip_memory2_1_s1_write                                   : out std_logic;                                        -- write
			onchip_memory2_1_s1_readdata                                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			onchip_memory2_1_s1_writedata                               : out std_logic_vector(31 downto 0);                    -- writedata
			onchip_memory2_1_s1_byteenable                              : out std_logic_vector(3 downto 0);                     -- byteenable
			onchip_memory2_1_s1_chipselect                              : out std_logic;                                        -- chipselect
			onchip_memory2_1_s1_clken                                   : out std_logic;                                        -- clken
			pin_s1_address                                              : out std_logic_vector(1 downto 0);                     -- address
			pin_s1_write                                                : out std_logic;                                        -- write
			pin_s1_readdata                                             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pin_s1_writedata                                            : out std_logic_vector(31 downto 0);                    -- writedata
			pin_s1_chipselect                                           : out std_logic;                                        -- chipselect
			pio_0_s1_address                                            : out std_logic_vector(1 downto 0);                     -- address
			pio_0_s1_write                                              : out std_logic;                                        -- write
			pio_0_s1_readdata                                           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pio_0_s1_writedata                                          : out std_logic_vector(31 downto 0);                    -- writedata
			pio_0_s1_chipselect                                         : out std_logic;                                        -- chipselect
			sysid_control_slave_address                                 : out std_logic_vector(0 downto 0);                     -- address
			sysid_control_slave_readdata                                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			timer_0_s1_address                                          : out std_logic_vector(2 downto 0);                     -- address
			timer_0_s1_write                                            : out std_logic;                                        -- write
			timer_0_s1_readdata                                         : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			timer_0_s1_writedata                                        : out std_logic_vector(15 downto 0);                    -- writedata
			timer_0_s1_chipselect                                       : out std_logic                                         -- chipselect
		);
	end component nios_system_mm_interconnect_0;

	component nios_system_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component nios_system_irq_mapper;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			reset_in1      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal sys_sdram_pll_0_sys_clk_clk                                                   : std_logic;                     -- sys_sdram_pll_0:sys_clk_clk -> [audio_0:clk, audio_and_video_config_0:clk, irq_mapper:clk, jtag_uart_0:clk, mm_interconnect_0:sys_sdram_pll_0_sys_clk_clk, new_sdram_controller_0:clk, nios2_gen2_0:clk, onchip_memory2_1:clk, pin:clk, pio_0:clk, rst_controller:clk, sysid:clock, timer_0:clk]
	signal nios2_gen2_0_data_master_readdata                                             : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	signal nios2_gen2_0_data_master_waitrequest                                          : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	signal nios2_gen2_0_data_master_debugaccess                                          : std_logic;                     -- nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	signal nios2_gen2_0_data_master_address                                              : std_logic_vector(26 downto 0); -- nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	signal nios2_gen2_0_data_master_byteenable                                           : std_logic_vector(3 downto 0);  -- nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	signal nios2_gen2_0_data_master_read                                                 : std_logic;                     -- nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	signal nios2_gen2_0_data_master_write                                                : std_logic;                     -- nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	signal nios2_gen2_0_data_master_writedata                                            : std_logic_vector(31 downto 0); -- nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	signal nios2_gen2_0_instruction_master_readdata                                      : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	signal nios2_gen2_0_instruction_master_waitrequest                                   : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	signal nios2_gen2_0_instruction_master_address                                       : std_logic_vector(26 downto 0); -- nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	signal nios2_gen2_0_instruction_master_read                                          : std_logic;                     -- nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	signal mm_interconnect_0_audio_0_avalon_audio_slave_chipselect                       : std_logic;                     -- mm_interconnect_0:audio_0_avalon_audio_slave_chipselect -> audio_0:chipselect
	signal mm_interconnect_0_audio_0_avalon_audio_slave_readdata                         : std_logic_vector(31 downto 0); -- audio_0:readdata -> mm_interconnect_0:audio_0_avalon_audio_slave_readdata
	signal mm_interconnect_0_audio_0_avalon_audio_slave_address                          : std_logic_vector(1 downto 0);  -- mm_interconnect_0:audio_0_avalon_audio_slave_address -> audio_0:address
	signal mm_interconnect_0_audio_0_avalon_audio_slave_read                             : std_logic;                     -- mm_interconnect_0:audio_0_avalon_audio_slave_read -> audio_0:read
	signal mm_interconnect_0_audio_0_avalon_audio_slave_write                            : std_logic;                     -- mm_interconnect_0:audio_0_avalon_audio_slave_write -> audio_0:write
	signal mm_interconnect_0_audio_0_avalon_audio_slave_writedata                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:audio_0_avalon_audio_slave_writedata -> audio_0:writedata
	signal mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_readdata    : std_logic_vector(31 downto 0); -- audio_and_video_config_0:readdata -> mm_interconnect_0:audio_and_video_config_0_avalon_av_config_slave_readdata
	signal mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_waitrequest : std_logic;                     -- audio_and_video_config_0:waitrequest -> mm_interconnect_0:audio_and_video_config_0_avalon_av_config_slave_waitrequest
	signal mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_address     : std_logic_vector(1 downto 0);  -- mm_interconnect_0:audio_and_video_config_0_avalon_av_config_slave_address -> audio_and_video_config_0:address
	signal mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_read        : std_logic;                     -- mm_interconnect_0:audio_and_video_config_0_avalon_av_config_slave_read -> audio_and_video_config_0:read
	signal mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_byteenable  : std_logic_vector(3 downto 0);  -- mm_interconnect_0:audio_and_video_config_0_avalon_av_config_slave_byteenable -> audio_and_video_config_0:byteenable
	signal mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_write       : std_logic;                     -- mm_interconnect_0:audio_and_video_config_0_avalon_av_config_slave_write -> audio_and_video_config_0:write
	signal mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_writedata   : std_logic_vector(31 downto 0); -- mm_interconnect_0:audio_and_video_config_0_avalon_av_config_slave_writedata -> audio_and_video_config_0:writedata
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect                    : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata                      : std_logic_vector(31 downto 0); -- jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest                   : std_logic;                     -- jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address                       : std_logic_vector(0 downto 0);  -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read                          : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write                         : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata                     : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	signal mm_interconnect_0_sysid_control_slave_readdata                                : std_logic_vector(31 downto 0); -- sysid:readdata -> mm_interconnect_0:sysid_control_slave_readdata
	signal mm_interconnect_0_sysid_control_slave_address                                 : std_logic_vector(0 downto 0);  -- mm_interconnect_0:sysid_control_slave_address -> sysid:address
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata                       : std_logic_vector(31 downto 0); -- nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest                    : std_logic;                     -- nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess                    : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address                        : std_logic_vector(8 downto 0);  -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read                           : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable                     : std_logic_vector(3 downto 0);  -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write                          : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata                      : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	signal mm_interconnect_0_onchip_memory2_1_s1_chipselect                              : std_logic;                     -- mm_interconnect_0:onchip_memory2_1_s1_chipselect -> onchip_memory2_1:chipselect
	signal mm_interconnect_0_onchip_memory2_1_s1_readdata                                : std_logic_vector(31 downto 0); -- onchip_memory2_1:readdata -> mm_interconnect_0:onchip_memory2_1_s1_readdata
	signal mm_interconnect_0_onchip_memory2_1_s1_address                                 : std_logic_vector(13 downto 0); -- mm_interconnect_0:onchip_memory2_1_s1_address -> onchip_memory2_1:address
	signal mm_interconnect_0_onchip_memory2_1_s1_byteenable                              : std_logic_vector(3 downto 0);  -- mm_interconnect_0:onchip_memory2_1_s1_byteenable -> onchip_memory2_1:byteenable
	signal mm_interconnect_0_onchip_memory2_1_s1_write                                   : std_logic;                     -- mm_interconnect_0:onchip_memory2_1_s1_write -> onchip_memory2_1:write
	signal mm_interconnect_0_onchip_memory2_1_s1_writedata                               : std_logic_vector(31 downto 0); -- mm_interconnect_0:onchip_memory2_1_s1_writedata -> onchip_memory2_1:writedata
	signal mm_interconnect_0_onchip_memory2_1_s1_clken                                   : std_logic;                     -- mm_interconnect_0:onchip_memory2_1_s1_clken -> onchip_memory2_1:clken
	signal mm_interconnect_0_pio_0_s1_chipselect                                         : std_logic;                     -- mm_interconnect_0:pio_0_s1_chipselect -> pio_0:chipselect
	signal mm_interconnect_0_pio_0_s1_readdata                                           : std_logic_vector(31 downto 0); -- pio_0:readdata -> mm_interconnect_0:pio_0_s1_readdata
	signal mm_interconnect_0_pio_0_s1_address                                            : std_logic_vector(1 downto 0);  -- mm_interconnect_0:pio_0_s1_address -> pio_0:address
	signal mm_interconnect_0_pio_0_s1_write                                              : std_logic;                     -- mm_interconnect_0:pio_0_s1_write -> mm_interconnect_0_pio_0_s1_write:in
	signal mm_interconnect_0_pio_0_s1_writedata                                          : std_logic_vector(31 downto 0); -- mm_interconnect_0:pio_0_s1_writedata -> pio_0:writedata
	signal mm_interconnect_0_new_sdram_controller_0_s1_chipselect                        : std_logic;                     -- mm_interconnect_0:new_sdram_controller_0_s1_chipselect -> new_sdram_controller_0:az_cs
	signal mm_interconnect_0_new_sdram_controller_0_s1_readdata                          : std_logic_vector(15 downto 0); -- new_sdram_controller_0:za_data -> mm_interconnect_0:new_sdram_controller_0_s1_readdata
	signal mm_interconnect_0_new_sdram_controller_0_s1_waitrequest                       : std_logic;                     -- new_sdram_controller_0:za_waitrequest -> mm_interconnect_0:new_sdram_controller_0_s1_waitrequest
	signal mm_interconnect_0_new_sdram_controller_0_s1_address                           : std_logic_vector(24 downto 0); -- mm_interconnect_0:new_sdram_controller_0_s1_address -> new_sdram_controller_0:az_addr
	signal mm_interconnect_0_new_sdram_controller_0_s1_read                              : std_logic;                     -- mm_interconnect_0:new_sdram_controller_0_s1_read -> mm_interconnect_0_new_sdram_controller_0_s1_read:in
	signal mm_interconnect_0_new_sdram_controller_0_s1_byteenable                        : std_logic_vector(1 downto 0);  -- mm_interconnect_0:new_sdram_controller_0_s1_byteenable -> mm_interconnect_0_new_sdram_controller_0_s1_byteenable:in
	signal mm_interconnect_0_new_sdram_controller_0_s1_readdatavalid                     : std_logic;                     -- new_sdram_controller_0:za_valid -> mm_interconnect_0:new_sdram_controller_0_s1_readdatavalid
	signal mm_interconnect_0_new_sdram_controller_0_s1_write                             : std_logic;                     -- mm_interconnect_0:new_sdram_controller_0_s1_write -> mm_interconnect_0_new_sdram_controller_0_s1_write:in
	signal mm_interconnect_0_new_sdram_controller_0_s1_writedata                         : std_logic_vector(15 downto 0); -- mm_interconnect_0:new_sdram_controller_0_s1_writedata -> new_sdram_controller_0:az_data
	signal mm_interconnect_0_timer_0_s1_chipselect                                       : std_logic;                     -- mm_interconnect_0:timer_0_s1_chipselect -> timer_0:chipselect
	signal mm_interconnect_0_timer_0_s1_readdata                                         : std_logic_vector(15 downto 0); -- timer_0:readdata -> mm_interconnect_0:timer_0_s1_readdata
	signal mm_interconnect_0_timer_0_s1_address                                          : std_logic_vector(2 downto 0);  -- mm_interconnect_0:timer_0_s1_address -> timer_0:address
	signal mm_interconnect_0_timer_0_s1_write                                            : std_logic;                     -- mm_interconnect_0:timer_0_s1_write -> mm_interconnect_0_timer_0_s1_write:in
	signal mm_interconnect_0_timer_0_s1_writedata                                        : std_logic_vector(15 downto 0); -- mm_interconnect_0:timer_0_s1_writedata -> timer_0:writedata
	signal mm_interconnect_0_pin_s1_chipselect                                           : std_logic;                     -- mm_interconnect_0:pin_s1_chipselect -> pin:chipselect
	signal mm_interconnect_0_pin_s1_readdata                                             : std_logic_vector(31 downto 0); -- pin:readdata -> mm_interconnect_0:pin_s1_readdata
	signal mm_interconnect_0_pin_s1_address                                              : std_logic_vector(1 downto 0);  -- mm_interconnect_0:pin_s1_address -> pin:address
	signal mm_interconnect_0_pin_s1_write                                                : std_logic;                     -- mm_interconnect_0:pin_s1_write -> mm_interconnect_0_pin_s1_write:in
	signal mm_interconnect_0_pin_s1_writedata                                            : std_logic_vector(31 downto 0); -- mm_interconnect_0:pin_s1_writedata -> pin:writedata
	signal irq_mapper_receiver0_irq                                                      : std_logic;                     -- jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                                      : std_logic;                     -- timer_0:irq -> irq_mapper:receiver1_irq
	signal nios2_gen2_0_irq_irq                                                          : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> nios2_gen2_0:irq
	signal rst_controller_reset_out_reset                                                : std_logic;                     -- rst_controller:reset_out -> [audio_0:reset, audio_and_video_config_0:reset, irq_mapper:reset, mm_interconnect_0:nios2_gen2_0_reset_reset_bridge_in_reset_reset, onchip_memory2_1:reset, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                                            : std_logic;                     -- rst_controller:reset_req -> [nios2_gen2_0:reset_req, onchip_memory2_1:reset_req, rst_translator:reset_req_in]
	signal nios2_gen2_0_debug_reset_request_reset                                        : std_logic;                     -- nios2_gen2_0:debug_reset_request -> rst_controller:reset_in0
	signal sys_sdram_pll_0_reset_source_reset                                            : std_logic;                     -- sys_sdram_pll_0:reset_source_reset -> rst_controller:reset_in1
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv                : std_logic;                     -- mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read:inv -> jtag_uart_0:av_read_n
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv               : std_logic;                     -- mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write:inv -> jtag_uart_0:av_write_n
	signal mm_interconnect_0_pio_0_s1_write_ports_inv                                    : std_logic;                     -- mm_interconnect_0_pio_0_s1_write:inv -> pio_0:write_n
	signal mm_interconnect_0_new_sdram_controller_0_s1_read_ports_inv                    : std_logic;                     -- mm_interconnect_0_new_sdram_controller_0_s1_read:inv -> new_sdram_controller_0:az_rd_n
	signal mm_interconnect_0_new_sdram_controller_0_s1_byteenable_ports_inv              : std_logic_vector(1 downto 0);  -- mm_interconnect_0_new_sdram_controller_0_s1_byteenable:inv -> new_sdram_controller_0:az_be_n
	signal mm_interconnect_0_new_sdram_controller_0_s1_write_ports_inv                   : std_logic;                     -- mm_interconnect_0_new_sdram_controller_0_s1_write:inv -> new_sdram_controller_0:az_wr_n
	signal mm_interconnect_0_timer_0_s1_write_ports_inv                                  : std_logic;                     -- mm_interconnect_0_timer_0_s1_write:inv -> timer_0:write_n
	signal mm_interconnect_0_pin_s1_write_ports_inv                                      : std_logic;                     -- mm_interconnect_0_pin_s1_write:inv -> pin:write_n
	signal rst_controller_reset_out_reset_ports_inv                                      : std_logic;                     -- rst_controller_reset_out_reset:inv -> [jtag_uart_0:rst_n, new_sdram_controller_0:reset_n, nios2_gen2_0:reset_n, pin:reset_n, pio_0:reset_n, sysid:reset_n, timer_0:reset_n]

begin

	audio_0 : component nios_system_audio_0
		port map (
			clk         => sys_sdram_pll_0_sys_clk_clk,                             --                clk.clk
			reset       => rst_controller_reset_out_reset,                          --              reset.reset
			address     => mm_interconnect_0_audio_0_avalon_audio_slave_address,    -- avalon_audio_slave.address
			chipselect  => mm_interconnect_0_audio_0_avalon_audio_slave_chipselect, --                   .chipselect
			read        => mm_interconnect_0_audio_0_avalon_audio_slave_read,       --                   .read
			write       => mm_interconnect_0_audio_0_avalon_audio_slave_write,      --                   .write
			writedata   => mm_interconnect_0_audio_0_avalon_audio_slave_writedata,  --                   .writedata
			readdata    => mm_interconnect_0_audio_0_avalon_audio_slave_readdata,   --                   .readdata
			irq         => open,                                                    --          interrupt.irq
			AUD_ADCDAT  => AUD_ADCDAT_to_the_audio_0,                               -- external_interface.export
			AUD_ADCLRCK => AUD_ADCLRCK_to_the_audio_0,                              --                   .export
			AUD_BCLK    => AUD_BCLK_to_the_audio_0,                                 --                   .export
			AUD_DACDAT  => AUD_DACDAT_from_the_audio_0,                             --                   .export
			AUD_DACLRCK => AUD_DACLRCK_to_the_audio_0                               --                   .export
		);

	audio_and_video_config_0 : component nios_system_audio_and_video_config_0
		port map (
			clk         => sys_sdram_pll_0_sys_clk_clk,                                                   --                    clk.clk
			reset       => rst_controller_reset_out_reset,                                                --                  reset.reset
			address     => mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_address,     -- avalon_av_config_slave.address
			byteenable  => mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_byteenable,  --                       .byteenable
			read        => mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_read,        --                       .read
			write       => mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_write,       --                       .write
			writedata   => mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_writedata,   --                       .writedata
			readdata    => mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_readdata,    --                       .readdata
			waitrequest => mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_waitrequest, --                       .waitrequest
			I2C_SDAT    => i2c_SDAT,                                                                      --     external_interface.export
			I2C_SCLK    => i2c_SCLK                                                                       --                       .export
		);

	jtag_uart_0 : component nios_system_jtag_uart_0
		port map (
			clk            => sys_sdram_pll_0_sys_clk_clk,                                     --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                        --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver0_irq                                         --               irq.irq
		);

	new_sdram_controller_0 : component nios_system_new_sdram_controller_0
		port map (
			clk            => sys_sdram_pll_0_sys_clk_clk,                                      --   clk.clk
			reset_n        => rst_controller_reset_out_reset_ports_inv,                         -- reset.reset_n
			az_addr        => mm_interconnect_0_new_sdram_controller_0_s1_address,              --    s1.address
			az_be_n        => mm_interconnect_0_new_sdram_controller_0_s1_byteenable_ports_inv, --      .byteenable_n
			az_cs          => mm_interconnect_0_new_sdram_controller_0_s1_chipselect,           --      .chipselect
			az_data        => mm_interconnect_0_new_sdram_controller_0_s1_writedata,            --      .writedata
			az_rd_n        => mm_interconnect_0_new_sdram_controller_0_s1_read_ports_inv,       --      .read_n
			az_wr_n        => mm_interconnect_0_new_sdram_controller_0_s1_write_ports_inv,      --      .write_n
			za_data        => mm_interconnect_0_new_sdram_controller_0_s1_readdata,             --      .readdata
			za_valid       => mm_interconnect_0_new_sdram_controller_0_s1_readdatavalid,        --      .readdatavalid
			za_waitrequest => mm_interconnect_0_new_sdram_controller_0_s1_waitrequest,          --      .waitrequest
			zs_addr        => sdram_addr,                                                       --  wire.export
			zs_ba          => sdram_ba,                                                         --      .export
			zs_cas_n       => sdram_cas_n,                                                      --      .export
			zs_cke         => sdram_cke,                                                        --      .export
			zs_cs_n        => sdram_cs_n,                                                       --      .export
			zs_dq          => sdram_dq,                                                         --      .export
			zs_dqm         => sdram_dqm,                                                        --      .export
			zs_ras_n       => sdram_ras_n,                                                      --      .export
			zs_we_n        => sdram_we_n                                                        --      .export
		);

	nios2_gen2_0 : component nios_system_nios2_gen2_0
		port map (
			clk                                 => sys_sdram_pll_0_sys_clk_clk,                                --                       clk.clk
			reset_n                             => rst_controller_reset_out_reset_ports_inv,                   --                     reset.reset_n
			reset_req                           => rst_controller_reset_out_reset_req,                         --                          .reset_req
			d_address                           => nios2_gen2_0_data_master_address,                           --               data_master.address
			d_byteenable                        => nios2_gen2_0_data_master_byteenable,                        --                          .byteenable
			d_read                              => nios2_gen2_0_data_master_read,                              --                          .read
			d_readdata                          => nios2_gen2_0_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => nios2_gen2_0_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => nios2_gen2_0_data_master_write,                             --                          .write
			d_writedata                         => nios2_gen2_0_data_master_writedata,                         --                          .writedata
			debug_mem_slave_debugaccess_to_roms => nios2_gen2_0_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => nios2_gen2_0_instruction_master_address,                    --        instruction_master.address
			i_read                              => nios2_gen2_0_instruction_master_read,                       --                          .read
			i_readdata                          => nios2_gen2_0_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => nios2_gen2_0_instruction_master_waitrequest,                --                          .waitrequest
			irq                                 => nios2_gen2_0_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => nios2_gen2_0_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                        -- custom_instruction_master.readra
		);

	onchip_memory2_1 : component nios_system_onchip_memory2_1
		port map (
			clk        => sys_sdram_pll_0_sys_clk_clk,                      --   clk1.clk
			address    => mm_interconnect_0_onchip_memory2_1_s1_address,    --     s1.address
			clken      => mm_interconnect_0_onchip_memory2_1_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_onchip_memory2_1_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_onchip_memory2_1_s1_write,      --       .write
			readdata   => mm_interconnect_0_onchip_memory2_1_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_onchip_memory2_1_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_onchip_memory2_1_s1_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,                   -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req,               --       .reset_req
			freeze     => '0'                                               -- (terminated)
		);

	pin : component nios_system_pin
		port map (
			clk        => sys_sdram_pll_0_sys_clk_clk,              --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address    => mm_interconnect_0_pin_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_pin_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_pin_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_pin_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_pin_s1_readdata,        --                    .readdata
			out_port   => pin_export                                -- external_connection.export
		);

	pio_0 : component nios_system_pio_0
		port map (
			clk        => sys_sdram_pll_0_sys_clk_clk,                --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,   --               reset.reset_n
			address    => mm_interconnect_0_pio_0_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_pio_0_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_pio_0_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_pio_0_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_pio_0_s1_readdata,        --                    .readdata
			in_port    => sw_export                                   -- external_connection.export
		);

	sys_sdram_pll_0 : component nios_system_sys_sdram_pll_0
		port map (
			ref_clk_clk        => clk_clk,                            --      ref_clk.clk
			ref_reset_reset    => reset_reset,                        --    ref_reset.reset
			sys_clk_clk        => sys_sdram_pll_0_sys_clk_clk,        --      sys_clk.clk
			sdram_clk_clk      => sdram_clk_clk,                      --    sdram_clk.clk
			reset_source_reset => sys_sdram_pll_0_reset_source_reset  -- reset_source.reset
		);

	sysid : component nios_system_sysid
		port map (
			clock    => sys_sdram_pll_0_sys_clk_clk,                      --           clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,         --         reset.reset_n
			readdata => mm_interconnect_0_sysid_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_0_sysid_control_slave_address(0)  --              .address
		);

	timer_0 : component nios_system_timer_0
		port map (
			clk        => sys_sdram_pll_0_sys_clk_clk,                  --   clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,     -- reset.reset_n
			address    => mm_interconnect_0_timer_0_s1_address,         --    s1.address
			writedata  => mm_interconnect_0_timer_0_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_0_timer_0_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_0_timer_0_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_0_timer_0_s1_write_ports_inv, --      .write_n
			irq        => irq_mapper_receiver1_irq                      --   irq.irq
		);

	mm_interconnect_0 : component nios_system_mm_interconnect_0
		port map (
			sys_sdram_pll_0_sys_clk_clk                                 => sys_sdram_pll_0_sys_clk_clk,                                                   --                         sys_sdram_pll_0_sys_clk.clk
			nios2_gen2_0_reset_reset_bridge_in_reset_reset              => rst_controller_reset_out_reset,                                                --        nios2_gen2_0_reset_reset_bridge_in_reset.reset
			nios2_gen2_0_data_master_address                            => nios2_gen2_0_data_master_address,                                              --                        nios2_gen2_0_data_master.address
			nios2_gen2_0_data_master_waitrequest                        => nios2_gen2_0_data_master_waitrequest,                                          --                                                .waitrequest
			nios2_gen2_0_data_master_byteenable                         => nios2_gen2_0_data_master_byteenable,                                           --                                                .byteenable
			nios2_gen2_0_data_master_read                               => nios2_gen2_0_data_master_read,                                                 --                                                .read
			nios2_gen2_0_data_master_readdata                           => nios2_gen2_0_data_master_readdata,                                             --                                                .readdata
			nios2_gen2_0_data_master_write                              => nios2_gen2_0_data_master_write,                                                --                                                .write
			nios2_gen2_0_data_master_writedata                          => nios2_gen2_0_data_master_writedata,                                            --                                                .writedata
			nios2_gen2_0_data_master_debugaccess                        => nios2_gen2_0_data_master_debugaccess,                                          --                                                .debugaccess
			nios2_gen2_0_instruction_master_address                     => nios2_gen2_0_instruction_master_address,                                       --                 nios2_gen2_0_instruction_master.address
			nios2_gen2_0_instruction_master_waitrequest                 => nios2_gen2_0_instruction_master_waitrequest,                                   --                                                .waitrequest
			nios2_gen2_0_instruction_master_read                        => nios2_gen2_0_instruction_master_read,                                          --                                                .read
			nios2_gen2_0_instruction_master_readdata                    => nios2_gen2_0_instruction_master_readdata,                                      --                                                .readdata
			audio_0_avalon_audio_slave_address                          => mm_interconnect_0_audio_0_avalon_audio_slave_address,                          --                      audio_0_avalon_audio_slave.address
			audio_0_avalon_audio_slave_write                            => mm_interconnect_0_audio_0_avalon_audio_slave_write,                            --                                                .write
			audio_0_avalon_audio_slave_read                             => mm_interconnect_0_audio_0_avalon_audio_slave_read,                             --                                                .read
			audio_0_avalon_audio_slave_readdata                         => mm_interconnect_0_audio_0_avalon_audio_slave_readdata,                         --                                                .readdata
			audio_0_avalon_audio_slave_writedata                        => mm_interconnect_0_audio_0_avalon_audio_slave_writedata,                        --                                                .writedata
			audio_0_avalon_audio_slave_chipselect                       => mm_interconnect_0_audio_0_avalon_audio_slave_chipselect,                       --                                                .chipselect
			audio_and_video_config_0_avalon_av_config_slave_address     => mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_address,     -- audio_and_video_config_0_avalon_av_config_slave.address
			audio_and_video_config_0_avalon_av_config_slave_write       => mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_write,       --                                                .write
			audio_and_video_config_0_avalon_av_config_slave_read        => mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_read,        --                                                .read
			audio_and_video_config_0_avalon_av_config_slave_readdata    => mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_readdata,    --                                                .readdata
			audio_and_video_config_0_avalon_av_config_slave_writedata   => mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_writedata,   --                                                .writedata
			audio_and_video_config_0_avalon_av_config_slave_byteenable  => mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_byteenable,  --                                                .byteenable
			audio_and_video_config_0_avalon_av_config_slave_waitrequest => mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_waitrequest, --                                                .waitrequest
			jtag_uart_0_avalon_jtag_slave_address                       => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address,                       --                   jtag_uart_0_avalon_jtag_slave.address
			jtag_uart_0_avalon_jtag_slave_write                         => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write,                         --                                                .write
			jtag_uart_0_avalon_jtag_slave_read                          => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read,                          --                                                .read
			jtag_uart_0_avalon_jtag_slave_readdata                      => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata,                      --                                                .readdata
			jtag_uart_0_avalon_jtag_slave_writedata                     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata,                     --                                                .writedata
			jtag_uart_0_avalon_jtag_slave_waitrequest                   => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest,                   --                                                .waitrequest
			jtag_uart_0_avalon_jtag_slave_chipselect                    => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect,                    --                                                .chipselect
			new_sdram_controller_0_s1_address                           => mm_interconnect_0_new_sdram_controller_0_s1_address,                           --                       new_sdram_controller_0_s1.address
			new_sdram_controller_0_s1_write                             => mm_interconnect_0_new_sdram_controller_0_s1_write,                             --                                                .write
			new_sdram_controller_0_s1_read                              => mm_interconnect_0_new_sdram_controller_0_s1_read,                              --                                                .read
			new_sdram_controller_0_s1_readdata                          => mm_interconnect_0_new_sdram_controller_0_s1_readdata,                          --                                                .readdata
			new_sdram_controller_0_s1_writedata                         => mm_interconnect_0_new_sdram_controller_0_s1_writedata,                         --                                                .writedata
			new_sdram_controller_0_s1_byteenable                        => mm_interconnect_0_new_sdram_controller_0_s1_byteenable,                        --                                                .byteenable
			new_sdram_controller_0_s1_readdatavalid                     => mm_interconnect_0_new_sdram_controller_0_s1_readdatavalid,                     --                                                .readdatavalid
			new_sdram_controller_0_s1_waitrequest                       => mm_interconnect_0_new_sdram_controller_0_s1_waitrequest,                       --                                                .waitrequest
			new_sdram_controller_0_s1_chipselect                        => mm_interconnect_0_new_sdram_controller_0_s1_chipselect,                        --                                                .chipselect
			nios2_gen2_0_debug_mem_slave_address                        => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address,                        --                    nios2_gen2_0_debug_mem_slave.address
			nios2_gen2_0_debug_mem_slave_write                          => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write,                          --                                                .write
			nios2_gen2_0_debug_mem_slave_read                           => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read,                           --                                                .read
			nios2_gen2_0_debug_mem_slave_readdata                       => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata,                       --                                                .readdata
			nios2_gen2_0_debug_mem_slave_writedata                      => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata,                      --                                                .writedata
			nios2_gen2_0_debug_mem_slave_byteenable                     => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable,                     --                                                .byteenable
			nios2_gen2_0_debug_mem_slave_waitrequest                    => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest,                    --                                                .waitrequest
			nios2_gen2_0_debug_mem_slave_debugaccess                    => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess,                    --                                                .debugaccess
			onchip_memory2_1_s1_address                                 => mm_interconnect_0_onchip_memory2_1_s1_address,                                 --                             onchip_memory2_1_s1.address
			onchip_memory2_1_s1_write                                   => mm_interconnect_0_onchip_memory2_1_s1_write,                                   --                                                .write
			onchip_memory2_1_s1_readdata                                => mm_interconnect_0_onchip_memory2_1_s1_readdata,                                --                                                .readdata
			onchip_memory2_1_s1_writedata                               => mm_interconnect_0_onchip_memory2_1_s1_writedata,                               --                                                .writedata
			onchip_memory2_1_s1_byteenable                              => mm_interconnect_0_onchip_memory2_1_s1_byteenable,                              --                                                .byteenable
			onchip_memory2_1_s1_chipselect                              => mm_interconnect_0_onchip_memory2_1_s1_chipselect,                              --                                                .chipselect
			onchip_memory2_1_s1_clken                                   => mm_interconnect_0_onchip_memory2_1_s1_clken,                                   --                                                .clken
			pin_s1_address                                              => mm_interconnect_0_pin_s1_address,                                              --                                          pin_s1.address
			pin_s1_write                                                => mm_interconnect_0_pin_s1_write,                                                --                                                .write
			pin_s1_readdata                                             => mm_interconnect_0_pin_s1_readdata,                                             --                                                .readdata
			pin_s1_writedata                                            => mm_interconnect_0_pin_s1_writedata,                                            --                                                .writedata
			pin_s1_chipselect                                           => mm_interconnect_0_pin_s1_chipselect,                                           --                                                .chipselect
			pio_0_s1_address                                            => mm_interconnect_0_pio_0_s1_address,                                            --                                        pio_0_s1.address
			pio_0_s1_write                                              => mm_interconnect_0_pio_0_s1_write,                                              --                                                .write
			pio_0_s1_readdata                                           => mm_interconnect_0_pio_0_s1_readdata,                                           --                                                .readdata
			pio_0_s1_writedata                                          => mm_interconnect_0_pio_0_s1_writedata,                                          --                                                .writedata
			pio_0_s1_chipselect                                         => mm_interconnect_0_pio_0_s1_chipselect,                                         --                                                .chipselect
			sysid_control_slave_address                                 => mm_interconnect_0_sysid_control_slave_address,                                 --                             sysid_control_slave.address
			sysid_control_slave_readdata                                => mm_interconnect_0_sysid_control_slave_readdata,                                --                                                .readdata
			timer_0_s1_address                                          => mm_interconnect_0_timer_0_s1_address,                                          --                                      timer_0_s1.address
			timer_0_s1_write                                            => mm_interconnect_0_timer_0_s1_write,                                            --                                                .write
			timer_0_s1_readdata                                         => mm_interconnect_0_timer_0_s1_readdata,                                         --                                                .readdata
			timer_0_s1_writedata                                        => mm_interconnect_0_timer_0_s1_writedata,                                        --                                                .writedata
			timer_0_s1_chipselect                                       => mm_interconnect_0_timer_0_s1_chipselect                                        --                                                .chipselect
		);

	irq_mapper : component nios_system_irq_mapper
		port map (
			clk           => sys_sdram_pll_0_sys_clk_clk,    --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,       -- receiver1.irq
			sender_irq    => nios2_gen2_0_irq_irq            --    sender.irq
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => nios2_gen2_0_debug_reset_request_reset, -- reset_in0.reset
			reset_in1      => sys_sdram_pll_0_reset_source_reset,     -- reset_in1.reset
			clk            => sys_sdram_pll_0_sys_clk_clk,            --       clk.clk
			reset_out      => rst_controller_reset_out_reset,         -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req,     --          .reset_req
			reset_req_in0  => '0',                                    -- (terminated)
			reset_req_in1  => '0',                                    -- (terminated)
			reset_in2      => '0',                                    -- (terminated)
			reset_req_in2  => '0',                                    -- (terminated)
			reset_in3      => '0',                                    -- (terminated)
			reset_req_in3  => '0',                                    -- (terminated)
			reset_in4      => '0',                                    -- (terminated)
			reset_req_in4  => '0',                                    -- (terminated)
			reset_in5      => '0',                                    -- (terminated)
			reset_req_in5  => '0',                                    -- (terminated)
			reset_in6      => '0',                                    -- (terminated)
			reset_req_in6  => '0',                                    -- (terminated)
			reset_in7      => '0',                                    -- (terminated)
			reset_req_in7  => '0',                                    -- (terminated)
			reset_in8      => '0',                                    -- (terminated)
			reset_req_in8  => '0',                                    -- (terminated)
			reset_in9      => '0',                                    -- (terminated)
			reset_req_in9  => '0',                                    -- (terminated)
			reset_in10     => '0',                                    -- (terminated)
			reset_req_in10 => '0',                                    -- (terminated)
			reset_in11     => '0',                                    -- (terminated)
			reset_req_in11 => '0',                                    -- (terminated)
			reset_in12     => '0',                                    -- (terminated)
			reset_req_in12 => '0',                                    -- (terminated)
			reset_in13     => '0',                                    -- (terminated)
			reset_req_in13 => '0',                                    -- (terminated)
			reset_in14     => '0',                                    -- (terminated)
			reset_req_in14 => '0',                                    -- (terminated)
			reset_in15     => '0',                                    -- (terminated)
			reset_req_in15 => '0'                                     -- (terminated)
		);

	mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;

	mm_interconnect_0_pio_0_s1_write_ports_inv <= not mm_interconnect_0_pio_0_s1_write;

	mm_interconnect_0_new_sdram_controller_0_s1_read_ports_inv <= not mm_interconnect_0_new_sdram_controller_0_s1_read;

	mm_interconnect_0_new_sdram_controller_0_s1_byteenable_ports_inv <= not mm_interconnect_0_new_sdram_controller_0_s1_byteenable;

	mm_interconnect_0_new_sdram_controller_0_s1_write_ports_inv <= not mm_interconnect_0_new_sdram_controller_0_s1_write;

	mm_interconnect_0_timer_0_s1_write_ports_inv <= not mm_interconnect_0_timer_0_s1_write;

	mm_interconnect_0_pin_s1_write_ports_inv <= not mm_interconnect_0_pin_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of nios_system
