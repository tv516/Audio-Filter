multiplier_inst : multiplier PORT MAP (
		dataa	 => dataa_sig,
		datab	 => datab_sig,
		result	 => result_sig
	);
